netcdf coordinate {
dimensions:
	Layer = 6 ;
variables:
	double Layer(Layer) ;
		Layer:long_name = "Layer Target Potential Density" ;
		Layer:units = "kg m-3" ;
		Layer:cartesian_axis = "Z" ;
		Layer:positive = "up" ;

// global attributes:
		:filename = "coordinate.nc" ;
data:

 Layer = 1025.5, 1027.1, 1027.5, 1027.8, 1028., 1028.2 ;
}
