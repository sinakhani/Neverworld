../NL_1deg/coordinate.cdl